library verilog;
use verilog.vl_types.all;
entity exp4_vlg_check_tst is
    port(
        bo              : in     vl_logic;
        df              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exp4_vlg_check_tst;
