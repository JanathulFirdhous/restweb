library verilog;
use verilog.vl_types.all;
entity exp2_vlg_check_tst is
    port(
        f1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exp2_vlg_check_tst;
