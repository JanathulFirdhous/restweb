library verilog;
use verilog.vl_types.all;
entity exp4_vlg_vec_tst is
end exp4_vlg_vec_tst;
