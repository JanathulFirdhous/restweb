library verilog;
use verilog.vl_types.all;
entity exp1_vlg_check_tst is
    port(
        f1              : in     vl_logic;
        f2              : in     vl_logic;
        f3              : in     vl_logic;
        f4              : in     vl_logic;
        f5              : in     vl_logic;
        f6              : in     vl_logic;
        f7              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end exp1_vlg_check_tst;
