library verilog;
use verilog.vl_types.all;
entity exp1_vlg_vec_tst is
end exp1_vlg_vec_tst;
